/* 
Verilog simulation of https://github.com/Johnlon/NESInterfaceAndPeripherals
*/
`ifndef V_GAMEPAD
`define V_GAMEPAD

`define EOF 32'hFFFF_FFFF 
`define NULL 0 
`define NL 10

`include "../lib/assertion.v"

`timescale 1ns/1ns

module gamepad_adapter #(parameter CONTROL_FILE="gamepad.control") (
    input  _OErandom, 
    input  _OEpad1, 
    input  _OEpad2, 
    output [7:0] Q
);

    function string strip;
        input string str;
    begin
        strip = str;
        if (str.len() > 0) begin
            if (str[str.len()-1] == `NL) begin
                strip = str.substr(0, str.len()-2); 
            end
        end
    end
    endfunction


    int fControl;
    int c, r;
    int tDelta;
    string strInput = "";
    string controlFile;
    integer iController;
    integer iControllerValue;
    reg [7:0] iController1Value;
    reg [7:0] iController2Value;
    localparam MAX_LINE_LENGTH=255;
    reg [8*MAX_LINE_LENGTH:0] line; /* Line of text read from file */ 


    initial 
    begin : file_block 
        if (! $value$plusargs("gamepad_control_file=%s", controlFile)) begin
            controlFile = CONTROL_FILE;
        end

        `ifndef verilator
                fControl = $fopenr(controlFile); 
        `endif


        if (fControl == `NULL) // If error opening file 
        begin
                $error("%9t ERROR ", $time, "failed opening file %s", controlFile);
                `FINISH_AND_RETURN(1);
                disable file_block; // Just quit 
        end

        while (fControl != `NULL)  
        begin
            c = $fgetc(fControl); 

            #100 // needed so that main loop gets a look in

            if (c != `EOF) 
            begin 
                if (c == "/") // identify controller  eg    c0=byte
                begin 
                    line="";
                    r = $fgets(line, fControl); 
                    strInput = strip(line);
                    $display("%9t ", $time, "GAMECONTROLLER: CONTROL RX: // %-s", strInput);
                end
                else if (c == "c") // identify controller  eg    c0=byte
                begin 
                    line="";
                    r = $fgets(line, fControl); 
                    strInput = strip(line);

                    r = $sscanf(strInput, "%1d=%02x", iController, iControllerValue);
                    if (r == 0) begin
                        $display("%9t ", $time, "GAMECONTROLLER: CONTROL RX: '%s' can't convert", strInput);
                    end

                    if (iController==1) begin
                        iController1Value = iControllerValue;
                        $display("%9t ", $time, "GAMECONTROLLER: CONTROL RX: 'c%s' :  controller 1 = %8b", strInput, iController1Value);
                    end
                    else if (iController==2) begin
                        iController2Value = iControllerValue;
                        $display("%9t ", $time, "GAMECONTROLLER: CONTROL RX: 'c%s' :  controller 2 = %8b", strInput, iController2Value);
                    end
                    else $display("%9t ", $time, "GAMECONTROLLER: CONTROL RX: 'c%s' :  %d is not a controller id", strInput, iController);


                end
                else if (c == "#") // sleep N ns
                begin
                    tDelta=0;
                    line="";
                    r = $fgets(line, fControl);  // consumes the line ending and space chars 
                    strInput = strip(line);

                    r = $sscanf(line,"%d\n", tDelta); 
                    #tDelta 
                    $display("%9t ", $time, "GAMECONTROLLER: CONTROL RX: '#%s' :  slept for %d", strInput, tDelta);
                    
                end
            end
        end
    end


    assign Q = _OEpad1 ? (_OEpad2 ? (_OErandom ? 8'bz: $random): iController2Value) : iController1Value;

endmodule

`endif

