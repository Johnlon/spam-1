
module main;
initial begin
$display("1");
$sleep(2999);
$display("2");
end
endmodule
