`include "exernal/ice-chips-verilog/Source-7400/74163.v"
`include "registerFile/syncRegisterFile.v"

`include "lib/assertion.v"

`timescale 1ns/100ps
`default_nettype none

module icarus_tb();
    
    
endmodule

