`include "hct74109.v" 
`include "../lib/assertion.v"
`timescale 1ns/1ns

module tb_jk;
   reg j;
   reg _k;
   reg clk=0;

   wire q, _q;
 
   // expected PD of device
   parameter PD=17;

    // must be longer than PD of device else malfunction
   parameter CLK_T=PD+1;

   parameter TEST_INTERVAL=CLK_T * 10;

   //always  #CLK_T clk = !clk;
    task clk_pulse;
    begin
        clk = 0;
        #CLK_T 
        clk = 1;
        #CLK_T 
        clk = 1; // repeat setting=1 otherwise syntax error cos can't have a delay as last item
    end
    endtask

 
   hct74109  jk0 ( .j(j),
                  ._k(_k),
                  .clk(clk),
                  .q(q),
                  ._q(_q)
    );
 
   initial begin
            // hold
      #TEST_INTERVAL 
        $display("hold mode");
        j <= 0;
        _k <= 1;

        clk_pulse();
        `Equals(q, 1'bx) // stays as X       
        clk_pulse();
        `Equals(q, 1'bx)
        clk_pulse();
        `Equals(q, 1'bx)
 
        // load reset Q=L
      #TEST_INTERVAL 
        $display("reset mode");
        j <= 0;
        _k <= 0;

        clk_pulse();
        `Equals(q, 1'b0)
        clk_pulse();
        `Equals(q, 1'b0)
        clk_pulse();
        `Equals(q, 1'b0)

        // load set Q=H
      #TEST_INTERVAL 
        $display("load mode");
        j <= 1;
        _k <= 1;

        clk_pulse();
        `Equals(q, 1'b1)
        clk_pulse();
        `Equals(q, 1'b1)
        clk_pulse();
        `Equals(q, 1'b1)

        // toggle
      #TEST_INTERVAL 
        $display("toggle mode");
        j <= 1;
        _k <= 0;

        `Equals(q, 1'b1)
        clk_pulse();
        `Equals(q, 1'b0)
        clk_pulse();
        `Equals(q, 1'b1)
        clk_pulse();
        `Equals(q, 1'b0)
        clk_pulse();
        `Equals(q, 1'b1)

      #TEST_INTERVAL $finish;
   end
 
   initial
      $monitor ($time, " clk ", clk, " j=%0d _k=%0d q=%0d", j, _k, q);

endmodule  
 

