// License: Mozilla Public License : Version 2.0
// Author : John Lonergan

module main;
initial begin
$display("1");
$sleep(2999);
$display("2");
end
endmodule
